
module not_gate(out,in);

    output [7:0] out;
    input [7:0] in;

    assign out = ~in;

endmodule





