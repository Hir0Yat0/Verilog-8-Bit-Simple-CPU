
module main (
    // ports

    

);
    
endmodule

