
module alu (
    // ports
    clk,
    alu_component_select,
    input_1,
    input_2,
    output_1,

);

    /* currently supports only add, multiply, and not add */    

    always @(posedge clk) begin
        
    end

    
endmodule







