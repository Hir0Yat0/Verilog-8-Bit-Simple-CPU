
// module decoder (
//     // ports
// );
    
// endmodule
