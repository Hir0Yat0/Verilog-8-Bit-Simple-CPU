
module or_gate(out,a,b); 

    output [7:0] out;
    input [7:0] a, b;

    assign out = a | b;

endmodule






