
module and_gate (
    // ports
    out,
    a,
    b,
);

    input a, b;
    output out;

    assign out = a & b;
    
endmodule
