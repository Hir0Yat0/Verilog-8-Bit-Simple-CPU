
module not_gate(out,in);

    output out;
    input in;

    assign out = ~in;

endmodule





