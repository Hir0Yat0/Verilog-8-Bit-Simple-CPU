
module alu (
    // ports
    // clk,
    alu_component_select,
    input_1,
    input_2,
    output_1,

);

    /* currently supports only add, multiply, and not add */    
    /* im pretty sure always @(*) check for any dependency inside blocks changes */
    always @(*) begin
        
    end

    
endmodule







